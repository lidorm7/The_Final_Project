Rom_X	Rom_X_inst (
	.address ( address_sig ),
	.clock ( clock_sig ),
	.q ( q_sig )
	);
